module audio_parallel_to_serial_testbench;
reg bck;
reg lrck;
reg  [15:0] datr;
reg  [15:0] datl;
wire out;
wire [3:0] temp;
wire temp2;
parameter stimDelay = 10;
audio_parallel_to_serial DUT(bck, lrck, out, datl, datr, temp,temp2);
initial
begin
//expected Rdata: 1100 1010 1100 1010
				 bck = 0; lrck = 0; datr=16'b1101010100101010; datl=16'b0000111100001111;
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; lrck=1;
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; lrck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1; datr=16'b0101010100101010; datl=16'b1000111100001111;
#(stimDelay) bck = 0; lrck = 1;
#(stimDelay) bck = 1; 
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 
#(stimDelay) bck = 1;
#(stimDelay) bck = 0; 

#100; //Let simulation finish
end

endmodule